module ALU(

    );
endmodule
